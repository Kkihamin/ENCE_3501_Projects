*** SPICE deck for cell ring_oscillator{sch} from library Lab6
*** Created on Sun Nov 05, 2023 22:25:08
*** Last revised on Fri Nov 10, 2023 12:01:44
*** Written on Fri Nov 10, 2023 12:11:17 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Lab6__NAND FROM CELL NAND{sch}
.SUBCKT Lab6__NAND A B Y
** GLOBAL 0
** GLOBAL vdd
Mnmos_2 Y A net_34 0 N_50n L=0.6U W=3U
Mnmos_3 net_34 B 0 0 N_50n L=0.6U W=3U
Mpmos_2 Y A vdd vdd P_50n L=0.6U W=3U
Mpmos_3 Y B vdd vdd P_50n L=0.6U W=3U
.ENDS Lab6__NAND

*** SUBCIRCUIT Lab6__NOT FROM CELL NOT{sch}
.SUBCKT Lab6__NOT A Y
** GLOBAL 0
** GLOBAL vdd
Mnmos_1 Y A 0 0 N_50n L=0.6U W=3U
Mpmos_1 Y A vdd vdd P_50n L=0.6U W=6U
.ENDS Lab6__NOT

.global 0 vdd

*** TOP LEVEL CELL: ring_oscillator{sch}
Cpoly2cap_0 0 net_0 10u
Cpoly2cap_1 0 net_31 10u
Cpoly2cap_2 0 net_35 10u
XNAND_0 osc En net_0 Lab6__NAND
XNOT_0 net_0 net_31 Lab6__NOT
XNOT_1 net_31 net_35 Lab6__NOT
XNOT_2 net_35 osc2 Lab6__NOT
XNOT_3 osc2 osc Lab6__NOT

* Spice Code nodes in cell cell 'ring_oscillator{sch}'
vdd vdd 0 dc 1
VEn En 0 dc 1
.tran 0 10
.include cmosedu_models.txt
.END
